
`include "alarm_trans.sv"
`include "alarm_gen.sv"
`include "alarm_intf.sv"
`include "alarm_bfm.sv"
`include "alarm_env.sv"
`include "alarm_test.sv"
`include "tb.sv"






